module RomNTT #(
parameter WIDTH_ADDR = 7,
parameter WIDTH_Data = 12
)(
input   logic   clk_i,
input   logic   rst_i,
input   logic   [WIDTH_ADDR - 1:0] address0,
input   logic   [WIDTH_ADDR - 1:0] address1,
input   logic   [WIDTH_ADDR - 1:0] address2,
input   logic   [WIDTH_ADDR - 1:0] address3,
input   logic   [WIDTH_ADDR - 1:0] address4,
input   logic   [WIDTH_ADDR - 1:0] address5,
input   logic   [WIDTH_ADDR - 1:0] address6,
input   logic   [WIDTH_ADDR - 1:0] address7,

output  logic   [WIDTH_Data - 1:0] q0,
output  logic   [WIDTH_Data - 1:0] q1,
output  logic   [WIDTH_Data - 1:0] q2,
output  logic   [WIDTH_Data - 1:0] q3,
output  logic   [WIDTH_Data - 1:0] q4,
output  logic   [WIDTH_Data - 1:0] q5,
output  logic   [WIDTH_Data - 1:0] q6,
output  logic   [WIDTH_Data - 1:0] q7
);

    logic [WIDTH_Data - 1:0] rom [0:127];

    always @(posedge clk_i) begin
        if(rst_i) begin
            rom[0] <= 12'd1;
            rom[1] <= 12'd1729;
            rom[2] <= 12'd2580;
            rom[3] <= 12'd3289;
            rom[4] <= 12'd2642;
            rom[5] <= 12'd630;
            rom[6] <= 12'd1897;
            rom[7] <= 12'd848;
            rom[8] <= 12'd1062;
            rom[9] <= 12'd1919;
            rom[10] <= 12'd193;
            rom[11] <= 12'd797;
            rom[12] <= 12'd2786;
            rom[13] <= 12'd3260;
            rom[14] <= 12'd569;
            rom[15] <= 12'd1746;
            rom[16] <= 12'd296;
            rom[17] <= 12'd2447;
            rom[18] <= 12'd1339;
            rom[19] <= 12'd1476;
            rom[20] <= 12'd3046;
            rom[21] <= 12'd56;
            rom[22] <= 12'd2240;
            rom[23] <= 12'd1333;
            rom[24] <= 12'd1426;
            rom[25] <= 12'd2094;
            rom[26] <= 12'd535;
            rom[27] <= 12'd2882;
            rom[28] <= 12'd2393;
            rom[29] <= 12'd2879;
            rom[30] <= 12'd1974;
            rom[31] <= 12'd821;
            rom[32] <= 12'd289;
            rom[33] <= 12'd331;
            rom[34] <= 12'd3253;
            rom[35] <= 12'd1756;
            rom[36] <= 12'd1197;
            rom[37] <= 12'd2304;
            rom[38] <= 12'd2277;
            rom[39] <= 12'd2055;
            rom[40] <= 12'd650;
            rom[41] <= 12'd1977;
            rom[42] <= 12'd2513;
            rom[43] <= 12'd632;
            rom[44] <= 12'd2865;
            rom[45] <= 12'd33;
            rom[46] <= 12'd1320;
            rom[47] <= 12'd1915;
            rom[48] <= 12'd2319;
            rom[49] <= 12'd1435;
            rom[50] <= 12'd807;
            rom[51] <= 12'd452;
            rom[52] <= 12'd1438;
            rom[53] <= 12'd2868;
            rom[54] <= 12'd1534;
            rom[55] <= 12'd2402;
            rom[56] <= 12'd2647;
            rom[57] <= 12'd2617;
            rom[58] <= 12'd1481;
            rom[59] <= 12'd648;
            rom[60] <= 12'd2474;
            rom[61] <= 12'd3110;
            rom[62] <= 12'd1227;
            rom[63] <= 12'd910;
            rom[64] <= 12'd17;
            rom[65] <= 12'd2761;
            rom[66] <= 12'd583;
            rom[67] <= 12'd2649;
            rom[68] <= 12'd1637;
            rom[69] <= 12'd723;
            rom[70] <= 12'd2288;
            rom[71] <= 12'd1100;
            rom[72] <= 12'd1409;
            rom[73] <= 12'd2662;
            rom[74] <= 12'd3281;
            rom[75] <= 12'd233;
            rom[76] <= 12'd756;
            rom[77] <= 12'd2156;
            rom[78] <= 12'd3015;
            rom[79] <= 12'd3050;
            rom[80] <= 12'd1703;
            rom[81] <= 12'd1651;
            rom[82] <= 12'd2789;
            rom[83] <= 12'd1789;
            rom[84] <= 12'd1847;
            rom[85] <= 12'd952;
            rom[86] <= 12'd1461;
            rom[87] <= 12'd2687;
            rom[88] <= 12'd939;
            rom[89] <= 12'd2308;
            rom[90] <= 12'd2437;
            rom[91] <= 12'd2388;
            rom[92] <= 12'd733;
            rom[93] <= 12'd2337;
            rom[94] <= 12'd268;
            rom[95] <= 12'd641;
            rom[96] <= 12'd1584;
            rom[97] <= 12'd2298;
            rom[98] <= 12'd2037;
            rom[99] <= 12'd3220;
            rom[100] <= 12'd375;
            rom[101] <= 12'd2549;
            rom[102] <= 12'd2090;
            rom[103] <= 12'd1645;
            rom[104] <= 12'd1063;
            rom[105] <= 12'd319;
            rom[106] <= 12'd2773;
            rom[107] <= 12'd757;
            rom[108] <= 12'd2099;
            rom[109] <= 12'd561;
            rom[110] <= 12'd2466;
            rom[111] <= 12'd2594;
            rom[112] <= 12'd2804;
            rom[113] <= 12'd1092;
            rom[114] <= 12'd403;
            rom[115] <= 12'd1026;
            rom[116] <= 12'd1143;
            rom[117] <= 12'd2150;
            rom[118] <= 12'd2775;
            rom[119] <= 12'd886;
            rom[120] <= 12'd1722;
            rom[121] <= 12'd1212;
            rom[122] <= 12'd1874;
            rom[123] <= 12'd1029;
            rom[124] <= 12'd2110;
            rom[125] <= 12'd2935;
            rom[126] <= 12'd885;
            rom[127] <= 12'd2154;
        end
    end
    // assign q = rom[address];
    assign q0 = rom[address0];
    assign q1 = rom[address1];
    assign q2 = rom[address2];
    assign q3 = rom[address3];
    assign q4 = rom[address4];
    assign q5 = rom[address5];
    assign q6 = rom[address6];
    assign q7 = rom[address7];
endmodule
