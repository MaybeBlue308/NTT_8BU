module BRAM_chain #(
    parameter DATA_WIDTH = 12,
    parameter INPUT_WIDTH = DATA_WIDTH * 16,
    parameter ADDR_WIDTH = 5,
    parameter DELAY_ADDR_WRITE = 7
    )(
    input logic                     clk_i,
    input logic                     rst_i,
    input logic [2:0]               mode_BRAM,
    input logic                     start_BRAM_chain,
    input logic                     start_BRAM_load,
    input logic                     start_BRAM_write,
    input logic                     we,
    input logic [DATA_WIDTH-1:0]    data_load_a,
    input logic [DATA_WIDTH-1:0]    data_load_b,
    input logic [ADDR_WIDTH-1:0]    addr_load_a,
    input logic [ADDR_WIDTH-1:0]    addr_load_b,
    /*--------------------------------*/
    input logic [ADDR_WIDTH-1:0]    data_in0, 
    input logic [ADDR_WIDTH-1:0]    data_in1, 
    input logic [ADDR_WIDTH-1:0]    data_in2,
    input logic [ADDR_WIDTH-1:0]    data_in3,
    input logic [ADDR_WIDTH-1:0]    data_in4,
    input logic [ADDR_WIDTH-1:0]    data_in5,
    input logic [ADDR_WIDTH-1:0]    data_in6,
    input logic [ADDR_WIDTH-1:0]    data_in7,
    input logic [ADDR_WIDTH-1:0]    data_in0B, 
    input logic [ADDR_WIDTH-1:0]    data_in1B, 
    input logic [ADDR_WIDTH-1:0]    data_in2B,
    input logic [ADDR_WIDTH-1:0]    data_in3B,
    input logic [ADDR_WIDTH-1:0]    data_in4B,
    input logic [ADDR_WIDTH-1:0]    data_in5B,
    input logic [ADDR_WIDTH-1:0]    data_in6B,
    input logic [ADDR_WIDTH-1:0]    data_in7B,
    /*--------------------------------*/
    input logic [ADDR_WIDTH-1:0]    addr_out0, 
    input logic [ADDR_WIDTH-1:0]    addr_out1, 
    input logic [ADDR_WIDTH-1:0]    addr_out2,
    input logic [ADDR_WIDTH-1:0]    addr_out3,
    input logic [ADDR_WIDTH-1:0]    addr_out4,
    input logic [ADDR_WIDTH-1:0]    addr_out5,
    input logic [ADDR_WIDTH-1:0]    addr_out6,
    input logic [ADDR_WIDTH-1:0]    addr_out7,
    input logic [ADDR_WIDTH-1:0]    addr_out0B, 
    input logic [ADDR_WIDTH-1:0]    addr_out1B, 
    input logic [ADDR_WIDTH-1:0]    addr_out2B,
    input logic [ADDR_WIDTH-1:0]    addr_out3B,
    input logic [ADDR_WIDTH-1:0]    addr_out4B,
    input logic [ADDR_WIDTH-1:0]    addr_out5B,
    input logic [ADDR_WIDTH-1:0]    addr_out6B,
    input logic [ADDR_WIDTH-1:0]    addr_out7B,    
    /*--------------------------------*/
    output logic [DATA_WIDTH-1:0]   data_bram0, 
    output logic [DATA_WIDTH-1:0]   data_bram1, 
    output logic [DATA_WIDTH-1:0]   data_bram2,
    output logic [DATA_WIDTH-1:0]   data_bram3, 
    output logic [DATA_WIDTH-1:0]   data_bram4, 
    output logic [DATA_WIDTH-1:0]   data_bram5, 
    output logic [DATA_WIDTH-1:0]   data_bram6,
    output logic [DATA_WIDTH-1:0]   data_bram7, 
    output logic [DATA_WIDTH-1:0]   data_bram0B, 
    output logic [DATA_WIDTH-1:0]   data_bram1B, 
    output logic [DATA_WIDTH-1:0]   data_bram2B,
    output logic [DATA_WIDTH-1:0]   data_bram3B,
    output logic [DATA_WIDTH-1:0]   data_bram4B,
    output logic [DATA_WIDTH-1:0]   data_bram5B,
    output logic [DATA_WIDTH-1:0]   data_bram6B,
    output logic [DATA_WIDTH-1:0]   data_bram7B,
    );

    logic [DATA_WIDTH]
    
    
endmodule